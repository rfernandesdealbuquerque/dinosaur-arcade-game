module LFSR_5bit(q7, q6, q5, q4, q3, clk, en, reset); //will vary bits 4 to 7 of output being 0000xxxx1111 - vary from 15 to 255

    input clk, en, reset;
    output q7, q6, q5, q4, q3;

    wire f;

    xnor XNOR(f, q7, q4);
    dffe_ref dff_7(.q(q7), .d(f), .clk(clk || reset), .en(1'b1), .clr(1'b0));
    dffe_ref dff_6(.q(q6), .d(q7), .clk(clk || reset), .en(1'b1), .clr(1'b0));
    dffe_ref dff_5(.q(q5), .d(q6), .clk(clk || reset), .en(1'b1), .clr(reset));
    dffe_ref dff_4(.q(q4), .d(q5), .clk(clk || reset), .en(1'b1), .clr(1'b0));
    dffe_ref dff_3(.q(q3), .d(q4), .clk(clk || reset), .en(1'b1), .clr(reset));


endmodule